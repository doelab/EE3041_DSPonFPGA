module IIR ();

endmodule
