module FIR ();

endmodule